library IEEE;
use IEEE.std_logic_1164.all;
entity Decompress is
    Port(clk: in std_logic;
        rst: in std_logic;
        din : in std_logic_vector(15 downto 0));
end entity Decompress;

architecture ArchIODecompress of Decompress is
begin
   
end ArchIODecompress;


