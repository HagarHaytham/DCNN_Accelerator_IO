library IEEE;
use IEEE.std_logic_1164.all;
entity IOInterface is
    Port(clk: in std_logic;
        rst: in std_logic;
        din : in std_logic_vector(15 downto 0));
end entity IOInterface;

architecture ArchIOInterface of IOInterface is
begin
   
end ArchIOInterface;


